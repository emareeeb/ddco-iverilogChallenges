module not2(y,a);
input a; output y;
assign y = ~ a;
endmodule 





